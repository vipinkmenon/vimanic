`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/04/2022 07:04:42 PM
// Design Name: 
// Module Name: angleLUT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module angleLUT #(parameter ampScale=1,stepSize=1,phase=0)(
input i_clk,
output [11:0] o_angle
);


reg[11:0] mem [0:1023];
reg [9:0] rdAddr;

assign o_angle = $signed($signed(mem[rdAddr])/$signed(ampScale));


always @(posedge i_clk)
begin
    if(rdAddr + stepSize > 1023)
        rdAddr <= 0;
    else
        rdAddr <= rdAddr + stepSize;
end

//LUT memory contains sine values in fixed
//point representation format.
//2 bit integer, 10 bit frac in 2's complement format 
//1024 samples for 2*pi radians  
initial
begin  
rdAddr = (1024*phase)/360;  
mem[0]= 0;
mem[1]= 12;
mem[2]= 25;
mem[3]= 37;
mem[4]= 50;
mem[5]= 62;
mem[6]= 75;
mem[7]= 87;
mem[8]= 100;
mem[9]= 113;
mem[10]= 125;
mem[11]= 138;
mem[12]= 150;
mem[13]= 163;
mem[14]= 175;
mem[15]= 188;
mem[16]= 200;
mem[17]= 213;
mem[18]= 225;
mem[19]= 238;
mem[20]= 250;
mem[21]= 263;
mem[22]= 275;
mem[23]= 288;
mem[24]= 300;
mem[25]= 312;
mem[26]= 325;
mem[27]= 337;
mem[28]= 350;
mem[29]= 362;
mem[30]= 374;
mem[31]= 387;
mem[32]= 399;
mem[33]= 411;
mem[34]= 424;
mem[35]= 436;
mem[36]= 448;
mem[37]= 460;
mem[38]= 473;
mem[39]= 485;
mem[40]= 497;
mem[41]= 509;
mem[42]= 521;
mem[43]= 534;
mem[44]= 546;
mem[45]= 558;
mem[46]= 570;
mem[47]= 582;
mem[48]= 594;
mem[49]= 606;
mem[50]= 618;
mem[51]= 630;
mem[52]= 642;
mem[53]= 654;
mem[54]= 666;
mem[55]= 678;
mem[56]= 689;
mem[57]= 701;
mem[58]= 713;
mem[59]= 725;
mem[60]= 737;
mem[61]= 748;
mem[62]= 760;
mem[63]= 772;
mem[64]= 783;
mem[65]= 795;
mem[66]= 806;
mem[67]= 818;
mem[68]= 829;
mem[69]= 841;
mem[70]= 852;
mem[71]= 864;
mem[72]= 875;
mem[73]= 886;
mem[74]= 898;
mem[75]= 909;
mem[76]= 920;
mem[77]= 932;
mem[78]= 943;
mem[79]= 954;
mem[80]= 965;
mem[81]= 976;
mem[82]= 987;
mem[83]= 998;
mem[84]= 1009;
mem[85]= 1020;
mem[86]= 1031;
mem[87]= 1042;
mem[88]= 1052;
mem[89]= 1063;
mem[90]= 1074;
mem[91]= 1085;
mem[92]= 1095;
mem[93]= 1106;
mem[94]= 1116;
mem[95]= 1127;
mem[96]= 1137;
mem[97]= 1148;
mem[98]= 1158;
mem[99]= 1168;
mem[100]= 1179;
mem[101]= 1189;
mem[102]= 1199;
mem[103]= 1209;
mem[104]= 1219;
mem[105]= 1230;
mem[106]= 1240;
mem[107]= 1250;
mem[108]= 1259;
mem[109]= 1269;
mem[110]= 1279;
mem[111]= 1289;
mem[112]= 1299;
mem[113]= 1308;
mem[114]= 1318;
mem[115]= 1328;
mem[116]= 1337;
mem[117]= 1347;
mem[118]= 1356;
mem[119]= 1366;
mem[120]= 1375;
mem[121]= 1384;
mem[122]= 1393;
mem[123]= 1403;
mem[124]= 1412;
mem[125]= 1421;
mem[126]= 1430;
mem[127]= 1439;
mem[128]= 1448;
mem[129]= 1457;
mem[130]= 1465;
mem[131]= 1474;
mem[132]= 1483;
mem[133]= 1491;
mem[134]= 1500;
mem[135]= 1509;
mem[136]= 1517;
mem[137]= 1525;
mem[138]= 1534;
mem[139]= 1542;
mem[140]= 1550;
mem[141]= 1558;
mem[142]= 1567;
mem[143]= 1575;
mem[144]= 1583;
mem[145]= 1591;
mem[146]= 1598;
mem[147]= 1606;
mem[148]= 1614;
mem[149]= 1622;
mem[150]= 1629;
mem[151]= 1637;
mem[152]= 1644;
mem[153]= 1652;
mem[154]= 1659;
mem[155]= 1667;
mem[156]= 1674;
mem[157]= 1681;
mem[158]= 1688;
mem[159]= 1695;
mem[160]= 1702;
mem[161]= 1709;
mem[162]= 1716;
mem[163]= 1723;
mem[164]= 1730;
mem[165]= 1736;
mem[166]= 1743;
mem[167]= 1750;
mem[168]= 1756;
mem[169]= 1763;
mem[170]= 1769;
mem[171]= 1775;
mem[172]= 1781;
mem[173]= 1788;
mem[174]= 1794;
mem[175]= 1800;
mem[176]= 1806;
mem[177]= 1812;
mem[178]= 1817;
mem[179]= 1823;
mem[180]= 1829;
mem[181]= 1834;
mem[182]= 1840;
mem[183]= 1845;
mem[184]= 1851;
mem[185]= 1856;
mem[186]= 1861;
mem[187]= 1867;
mem[188]= 1872;
mem[189]= 1877;
mem[190]= 1882;
mem[191]= 1887;
mem[192]= 1892;
mem[193]= 1896;
mem[194]= 1901;
mem[195]= 1906;
mem[196]= 1910;
mem[197]= 1915;
mem[198]= 1919;
mem[199]= 1924;
mem[200]= 1928;
mem[201]= 1932;
mem[202]= 1936;
mem[203]= 1940;
mem[204]= 1944;
mem[205]= 1948;
mem[206]= 1952;
mem[207]= 1956;
mem[208]= 1959;
mem[209]= 1963;
mem[210]= 1966;
mem[211]= 1970;
mem[212]= 1973;
mem[213]= 1977;
mem[214]= 1980;
mem[215]= 1983;
mem[216]= 1986;
mem[217]= 1989;
mem[218]= 1992;
mem[219]= 1995;
mem[220]= 1998;
mem[221]= 2000;
mem[222]= 2003;
mem[223]= 2006;
mem[224]= 2008;
mem[225]= 2011;
mem[226]= 2013;
mem[227]= 2015;
mem[228]= 2017;
mem[229]= 2019;
mem[230]= 2021;
mem[231]= 2023;
mem[232]= 2025;
mem[233]= 2027;
mem[234]= 2029;
mem[235]= 2031;
mem[236]= 2032;
mem[237]= 2034;
mem[238]= 2035;
mem[239]= 2036;
mem[240]= 2038;
mem[241]= 2039;
mem[242]= 2040;
mem[243]= 2041;
mem[244]= 2042;
mem[245]= 2043;
mem[246]= 2044;
mem[247]= 2044;
mem[248]= 2045;
mem[249]= 2046;
mem[250]= 2046;
mem[251]= 2047;
mem[252]= 2047;
mem[253]= 2047;
mem[254]= 2047;
mem[255]= 2047;
mem[256]= 2047;
mem[257]= 2047;
mem[258]= 2047;
mem[259]= 2047;
mem[260]= 2047;
mem[261]= 2047;
mem[262]= 2046;
mem[263]= 2046;
mem[264]= 2045;
mem[265]= 2044;
mem[266]= 2044;
mem[267]= 2043;
mem[268]= 2042;
mem[269]= 2041;
mem[270]= 2040;
mem[271]= 2039;
mem[272]= 2038;
mem[273]= 2036;
mem[274]= 2035;
mem[275]= 2034;
mem[276]= 2032;
mem[277]= 2031;
mem[278]= 2029;
mem[279]= 2027;
mem[280]= 2025;
mem[281]= 2023;
mem[282]= 2021;
mem[283]= 2019;
mem[284]= 2017;
mem[285]= 2015;
mem[286]= 2013;
mem[287]= 2011;
mem[288]= 2008;
mem[289]= 2006;
mem[290]= 2003;
mem[291]= 2000;
mem[292]= 1998;
mem[293]= 1995;
mem[294]= 1992;
mem[295]= 1989;
mem[296]= 1986;
mem[297]= 1983;
mem[298]= 1980;
mem[299]= 1977;
mem[300]= 1973;
mem[301]= 1970;
mem[302]= 1966;
mem[303]= 1963;
mem[304]= 1959;
mem[305]= 1956;
mem[306]= 1952;
mem[307]= 1948;
mem[308]= 1944;
mem[309]= 1940;
mem[310]= 1936;
mem[311]= 1932;
mem[312]= 1928;
mem[313]= 1924;
mem[314]= 1919;
mem[315]= 1915;
mem[316]= 1910;
mem[317]= 1906;
mem[318]= 1901;
mem[319]= 1896;
mem[320]= 1892;
mem[321]= 1887;
mem[322]= 1882;
mem[323]= 1877;
mem[324]= 1872;
mem[325]= 1867;
mem[326]= 1861;
mem[327]= 1856;
mem[328]= 1851;
mem[329]= 1845;
mem[330]= 1840;
mem[331]= 1834;
mem[332]= 1829;
mem[333]= 1823;
mem[334]= 1817;
mem[335]= 1812;
mem[336]= 1806;
mem[337]= 1800;
mem[338]= 1794;
mem[339]= 1788;
mem[340]= 1781;
mem[341]= 1775;
mem[342]= 1769;
mem[343]= 1763;
mem[344]= 1756;
mem[345]= 1750;
mem[346]= 1743;
mem[347]= 1736;
mem[348]= 1730;
mem[349]= 1723;
mem[350]= 1716;
mem[351]= 1709;
mem[352]= 1702;
mem[353]= 1695;
mem[354]= 1688;
mem[355]= 1681;
mem[356]= 1674;
mem[357]= 1667;
mem[358]= 1659;
mem[359]= 1652;
mem[360]= 1644;
mem[361]= 1637;
mem[362]= 1629;
mem[363]= 1622;
mem[364]= 1614;
mem[365]= 1606;
mem[366]= 1598;
mem[367]= 1591;
mem[368]= 1583;
mem[369]= 1575;
mem[370]= 1567;
mem[371]= 1558;
mem[372]= 1550;
mem[373]= 1542;
mem[374]= 1534;
mem[375]= 1525;
mem[376]= 1517;
mem[377]= 1509;
mem[378]= 1500;
mem[379]= 1491;
mem[380]= 1483;
mem[381]= 1474;
mem[382]= 1465;
mem[383]= 1457;
mem[384]= 1448;
mem[385]= 1439;
mem[386]= 1430;
mem[387]= 1421;
mem[388]= 1412;
mem[389]= 1403;
mem[390]= 1393;
mem[391]= 1384;
mem[392]= 1375;
mem[393]= 1366;
mem[394]= 1356;
mem[395]= 1347;
mem[396]= 1337;
mem[397]= 1328;
mem[398]= 1318;
mem[399]= 1308;
mem[400]= 1299;
mem[401]= 1289;
mem[402]= 1279;
mem[403]= 1269;
mem[404]= 1259;
mem[405]= 1250;
mem[406]= 1240;
mem[407]= 1230;
mem[408]= 1219;
mem[409]= 1209;
mem[410]= 1199;
mem[411]= 1189;
mem[412]= 1179;
mem[413]= 1168;
mem[414]= 1158;
mem[415]= 1148;
mem[416]= 1137;
mem[417]= 1127;
mem[418]= 1116;
mem[419]= 1106;
mem[420]= 1095;
mem[421]= 1085;
mem[422]= 1074;
mem[423]= 1063;
mem[424]= 1052;
mem[425]= 1042;
mem[426]= 1031;
mem[427]= 1020;
mem[428]= 1009;
mem[429]= 998;
mem[430]= 987;
mem[431]= 976;
mem[432]= 965;
mem[433]= 954;
mem[434]= 943;
mem[435]= 932;
mem[436]= 920;
mem[437]= 909;
mem[438]= 898;
mem[439]= 886;
mem[440]= 875;
mem[441]= 864;
mem[442]= 852;
mem[443]= 841;
mem[444]= 829;
mem[445]= 818;
mem[446]= 806;
mem[447]= 795;
mem[448]= 783;
mem[449]= 772;
mem[450]= 760;
mem[451]= 748;
mem[452]= 737;
mem[453]= 725;
mem[454]= 713;
mem[455]= 701;
mem[456]= 689;
mem[457]= 678;
mem[458]= 666;
mem[459]= 654;
mem[460]= 642;
mem[461]= 630;
mem[462]= 618;
mem[463]= 606;
mem[464]= 594;
mem[465]= 582;
mem[466]= 570;
mem[467]= 558;
mem[468]= 546;
mem[469]= 534;
mem[470]= 521;
mem[471]= 509;
mem[472]= 497;
mem[473]= 485;
mem[474]= 473;
mem[475]= 460;
mem[476]= 448;
mem[477]= 436;
mem[478]= 424;
mem[479]= 411;
mem[480]= 399;
mem[481]= 387;
mem[482]= 374;
mem[483]= 362;
mem[484]= 350;
mem[485]= 337;
mem[486]= 325;
mem[487]= 312;
mem[488]= 300;
mem[489]= 288;
mem[490]= 275;
mem[491]= 263;
mem[492]= 250;
mem[493]= 238;
mem[494]= 225;
mem[495]= 213;
mem[496]= 200;
mem[497]= 188;
mem[498]= 175;
mem[499]= 163;
mem[500]= 150;
mem[501]= 138;
mem[502]= 125;
mem[503]= 113;
mem[504]= 100;
mem[505]= 87;
mem[506]= 75;
mem[507]= 62;
mem[508]= 50;
mem[509]= 37;
mem[510]= 25;
mem[511]= 12;
mem[512]= 0;
mem[513]= 4084;
mem[514]= 4071;
mem[515]= 4059;
mem[516]= 4046;
mem[517]= 4034;
mem[518]= 4021;
mem[519]= 4009;
mem[520]= 3996;
mem[521]= 3983;
mem[522]= 3971;
mem[523]= 3958;
mem[524]= 3946;
mem[525]= 3933;
mem[526]= 3921;
mem[527]= 3908;
mem[528]= 3896;
mem[529]= 3883;
mem[530]= 3871;
mem[531]= 3858;
mem[532]= 3846;
mem[533]= 3833;
mem[534]= 3821;
mem[535]= 3808;
mem[536]= 3796;
mem[537]= 3784;
mem[538]= 3771;
mem[539]= 3759;
mem[540]= 3746;
mem[541]= 3734;
mem[542]= 3722;
mem[543]= 3709;
mem[544]= 3697;
mem[545]= 3685;
mem[546]= 3672;
mem[547]= 3660;
mem[548]= 3648;
mem[549]= 3636;
mem[550]= 3623;
mem[551]= 3611;
mem[552]= 3599;
mem[553]= 3587;
mem[554]= 3575;
mem[555]= 3562;
mem[556]= 3550;
mem[557]= 3538;
mem[558]= 3526;
mem[559]= 3514;
mem[560]= 3502;
mem[561]= 3490;
mem[562]= 3478;
mem[563]= 3466;
mem[564]= 3454;
mem[565]= 3442;
mem[566]= 3430;
mem[567]= 3418;
mem[568]= 3407;
mem[569]= 3395;
mem[570]= 3383;
mem[571]= 3371;
mem[572]= 3359;
mem[573]= 3348;
mem[574]= 3336;
mem[575]= 3324;
mem[576]= 3313;
mem[577]= 3301;
mem[578]= 3290;
mem[579]= 3278;
mem[580]= 3267;
mem[581]= 3255;
mem[582]= 3244;
mem[583]= 3232;
mem[584]= 3221;
mem[585]= 3210;
mem[586]= 3198;
mem[587]= 3187;
mem[588]= 3176;
mem[589]= 3164;
mem[590]= 3153;
mem[591]= 3142;
mem[592]= 3131;
mem[593]= 3120;
mem[594]= 3109;
mem[595]= 3098;
mem[596]= 3087;
mem[597]= 3076;
mem[598]= 3065;
mem[599]= 3054;
mem[600]= 3044;
mem[601]= 3033;
mem[602]= 3022;
mem[603]= 3011;
mem[604]= 3001;
mem[605]= 2990;
mem[606]= 2980;
mem[607]= 2969;
mem[608]= 2959;
mem[609]= 2948;
mem[610]= 2938;
mem[611]= 2928;
mem[612]= 2917;
mem[613]= 2907;
mem[614]= 2897;
mem[615]= 2887;
mem[616]= 2877;
mem[617]= 2866;
mem[618]= 2856;
mem[619]= 2846;
mem[620]= 2837;
mem[621]= 2827;
mem[622]= 2817;
mem[623]= 2807;
mem[624]= 2797;
mem[625]= 2788;
mem[626]= 2778;
mem[627]= 2768;
mem[628]= 2759;
mem[629]= 2749;
mem[630]= 2740;
mem[631]= 2730;
mem[632]= 2721;
mem[633]= 2712;
mem[634]= 2703;
mem[635]= 2693;
mem[636]= 2684;
mem[637]= 2675;
mem[638]= 2666;
mem[639]= 2657;
mem[640]= 2648;
mem[641]= 2639;
mem[642]= 2631;
mem[643]= 2622;
mem[644]= 2613;
mem[645]= 2605;
mem[646]= 2596;
mem[647]= 2587;
mem[648]= 2579;
mem[649]= 2571;
mem[650]= 2562;
mem[651]= 2554;
mem[652]= 2546;
mem[653]= 2538;
mem[654]= 2529;
mem[655]= 2521;
mem[656]= 2513;
mem[657]= 2505;
mem[658]= 2498;
mem[659]= 2490;
mem[660]= 2482;
mem[661]= 2474;
mem[662]= 2467;
mem[663]= 2459;
mem[664]= 2452;
mem[665]= 2444;
mem[666]= 2437;
mem[667]= 2429;
mem[668]= 2422;
mem[669]= 2415;
mem[670]= 2408;
mem[671]= 2401;
mem[672]= 2394;
mem[673]= 2387;
mem[674]= 2380;
mem[675]= 2373;
mem[676]= 2366;
mem[677]= 2360;
mem[678]= 2353;
mem[679]= 2346;
mem[680]= 2340;
mem[681]= 2333;
mem[682]= 2327;
mem[683]= 2321;
mem[684]= 2315;
mem[685]= 2308;
mem[686]= 2302;
mem[687]= 2296;
mem[688]= 2290;
mem[689]= 2284;
mem[690]= 2279;
mem[691]= 2273;
mem[692]= 2267;
mem[693]= 2262;
mem[694]= 2256;
mem[695]= 2251;
mem[696]= 2245;
mem[697]= 2240;
mem[698]= 2235;
mem[699]= 2229;
mem[700]= 2224;
mem[701]= 2219;
mem[702]= 2214;
mem[703]= 2209;
mem[704]= 2204;
mem[705]= 2200;
mem[706]= 2195;
mem[707]= 2190;
mem[708]= 2186;
mem[709]= 2181;
mem[710]= 2177;
mem[711]= 2172;
mem[712]= 2168;
mem[713]= 2164;
mem[714]= 2160;
mem[715]= 2156;
mem[716]= 2152;
mem[717]= 2148;
mem[718]= 2144;
mem[719]= 2140;
mem[720]= 2137;
mem[721]= 2133;
mem[722]= 2130;
mem[723]= 2126;
mem[724]= 2123;
mem[725]= 2119;
mem[726]= 2116;
mem[727]= 2113;
mem[728]= 2110;
mem[729]= 2107;
mem[730]= 2104;
mem[731]= 2101;
mem[732]= 2098;
mem[733]= 2096;
mem[734]= 2093;
mem[735]= 2090;
mem[736]= 2088;
mem[737]= 2085;
mem[738]= 2083;
mem[739]= 2081;
mem[740]= 2079;
mem[741]= 2077;
mem[742]= 2075;
mem[743]= 2073;
mem[744]= 2071;
mem[745]= 2069;
mem[746]= 2067;
mem[747]= 2065;
mem[748]= 2064;
mem[749]= 2062;
mem[750]= 2061;
mem[751]= 2060;
mem[752]= 2058;
mem[753]= 2057;
mem[754]= 2056;
mem[755]= 2055;
mem[756]= 2054;
mem[757]= 2053;
mem[758]= 2052;
mem[759]= 2052;
mem[760]= 2051;
mem[761]= 2050;
mem[762]= 2050;
mem[763]= 2049;
mem[764]= 2049;
mem[765]= 2049;
mem[766]= 2049;
mem[767]= 2049;
mem[768]= 2048;
mem[769]= 2049;
mem[770]= 2049;
mem[771]= 2049;
mem[772]= 2049;
mem[773]= 2049;
mem[774]= 2050;
mem[775]= 2050;
mem[776]= 2051;
mem[777]= 2052;
mem[778]= 2052;
mem[779]= 2053;
mem[780]= 2054;
mem[781]= 2055;
mem[782]= 2056;
mem[783]= 2057;
mem[784]= 2058;
mem[785]= 2060;
mem[786]= 2061;
mem[787]= 2062;
mem[788]= 2064;
mem[789]= 2065;
mem[790]= 2067;
mem[791]= 2069;
mem[792]= 2071;
mem[793]= 2073;
mem[794]= 2075;
mem[795]= 2077;
mem[796]= 2079;
mem[797]= 2081;
mem[798]= 2083;
mem[799]= 2085;
mem[800]= 2088;
mem[801]= 2090;
mem[802]= 2093;
mem[803]= 2096;
mem[804]= 2098;
mem[805]= 2101;
mem[806]= 2104;
mem[807]= 2107;
mem[808]= 2110;
mem[809]= 2113;
mem[810]= 2116;
mem[811]= 2119;
mem[812]= 2123;
mem[813]= 2126;
mem[814]= 2130;
mem[815]= 2133;
mem[816]= 2137;
mem[817]= 2140;
mem[818]= 2144;
mem[819]= 2148;
mem[820]= 2152;
mem[821]= 2156;
mem[822]= 2160;
mem[823]= 2164;
mem[824]= 2168;
mem[825]= 2172;
mem[826]= 2177;
mem[827]= 2181;
mem[828]= 2186;
mem[829]= 2190;
mem[830]= 2195;
mem[831]= 2200;
mem[832]= 2204;
mem[833]= 2209;
mem[834]= 2214;
mem[835]= 2219;
mem[836]= 2224;
mem[837]= 2229;
mem[838]= 2235;
mem[839]= 2240;
mem[840]= 2245;
mem[841]= 2251;
mem[842]= 2256;
mem[843]= 2262;
mem[844]= 2267;
mem[845]= 2273;
mem[846]= 2279;
mem[847]= 2284;
mem[848]= 2290;
mem[849]= 2296;
mem[850]= 2302;
mem[851]= 2308;
mem[852]= 2315;
mem[853]= 2321;
mem[854]= 2327;
mem[855]= 2333;
mem[856]= 2340;
mem[857]= 2346;
mem[858]= 2353;
mem[859]= 2360;
mem[860]= 2366;
mem[861]= 2373;
mem[862]= 2380;
mem[863]= 2387;
mem[864]= 2394;
mem[865]= 2401;
mem[866]= 2408;
mem[867]= 2415;
mem[868]= 2422;
mem[869]= 2429;
mem[870]= 2437;
mem[871]= 2444;
mem[872]= 2452;
mem[873]= 2459;
mem[874]= 2467;
mem[875]= 2474;
mem[876]= 2482;
mem[877]= 2490;
mem[878]= 2498;
mem[879]= 2505;
mem[880]= 2513;
mem[881]= 2521;
mem[882]= 2529;
mem[883]= 2538;
mem[884]= 2546;
mem[885]= 2554;
mem[886]= 2562;
mem[887]= 2571;
mem[888]= 2579;
mem[889]= 2587;
mem[890]= 2596;
mem[891]= 2605;
mem[892]= 2613;
mem[893]= 2622;
mem[894]= 2631;
mem[895]= 2639;
mem[896]= 2648;
mem[897]= 2657;
mem[898]= 2666;
mem[899]= 2675;
mem[900]= 2684;
mem[901]= 2693;
mem[902]= 2703;
mem[903]= 2712;
mem[904]= 2721;
mem[905]= 2730;
mem[906]= 2740;
mem[907]= 2749;
mem[908]= 2759;
mem[909]= 2768;
mem[910]= 2778;
mem[911]= 2788;
mem[912]= 2797;
mem[913]= 2807;
mem[914]= 2817;
mem[915]= 2827;
mem[916]= 2837;
mem[917]= 2846;
mem[918]= 2856;
mem[919]= 2866;
mem[920]= 2877;
mem[921]= 2887;
mem[922]= 2897;
mem[923]= 2907;
mem[924]= 2917;
mem[925]= 2928;
mem[926]= 2938;
mem[927]= 2948;
mem[928]= 2959;
mem[929]= 2969;
mem[930]= 2980;
mem[931]= 2990;
mem[932]= 3001;
mem[933]= 3011;
mem[934]= 3022;
mem[935]= 3033;
mem[936]= 3044;
mem[937]= 3054;
mem[938]= 3065;
mem[939]= 3076;
mem[940]= 3087;
mem[941]= 3098;
mem[942]= 3109;
mem[943]= 3120;
mem[944]= 3131;
mem[945]= 3142;
mem[946]= 3153;
mem[947]= 3164;
mem[948]= 3176;
mem[949]= 3187;
mem[950]= 3198;
mem[951]= 3210;
mem[952]= 3221;
mem[953]= 3232;
mem[954]= 3244;
mem[955]= 3255;
mem[956]= 3267;
mem[957]= 3278;
mem[958]= 3290;
mem[959]= 3301;
mem[960]= 3313;
mem[961]= 3324;
mem[962]= 3336;
mem[963]= 3348;
mem[964]= 3359;
mem[965]= 3371;
mem[966]= 3383;
mem[967]= 3395;
mem[968]= 3407;
mem[969]= 3418;
mem[970]= 3430;
mem[971]= 3442;
mem[972]= 3454;
mem[973]= 3466;
mem[974]= 3478;
mem[975]= 3490;
mem[976]= 3502;
mem[977]= 3514;
mem[978]= 3526;
mem[979]= 3538;
mem[980]= 3550;
mem[981]= 3562;
mem[982]= 3575;
mem[983]= 3587;
mem[984]= 3599;
mem[985]= 3611;
mem[986]= 3623;
mem[987]= 3636;
mem[988]= 3648;
mem[989]= 3660;
mem[990]= 3672;
mem[991]= 3685;
mem[992]= 3697;
mem[993]= 3709;
mem[994]= 3722;
mem[995]= 3734;
mem[996]= 3746;
mem[997]= 3759;
mem[998]= 3771;
mem[999]= 3784;
mem[1000]= 3796;
mem[1001]= 3808;
mem[1002]= 3821;
mem[1003]= 3833;
mem[1004]= 3846;
mem[1005]= 3858;
mem[1006]= 3871;
mem[1007]= 3883;
mem[1008]= 3896;
mem[1009]= 3908;
mem[1010]= 3921;
mem[1011]= 3933;
mem[1012]= 3946;
mem[1013]= 3958;
mem[1014]= 3971;
mem[1015]= 3983;
mem[1016]= 3996;
mem[1017]= 4009;
mem[1018]= 4021;
mem[1019]= 4034;
mem[1020]= 4046;
mem[1021]= 4059;
mem[1022]= 4071;
mem[1023]= 4084;
end
    
    
    
endmodule